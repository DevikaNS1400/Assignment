`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mux_4_1(
output Y,
input S1,S0,I3,I2,I1,I0
    );
assign Y=(S1)?((S0)?I3:I2):((S0)?I1:I0);
endmodule
