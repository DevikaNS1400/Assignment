`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
//////////////////////////////////////////////////////////////////////////////////


module mod_N_comp #(parameter N=4)(
output aeb,alb,agb,
input [N-1:0]a,b
 );
 assign aeb=((a<=b)&&(a>=b))?1'b1:0;
 assign alb=(a<b)?1'b1:0;
 assign agb=(a>=b)?1'b1:0; 
endmodule
