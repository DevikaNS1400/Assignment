`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_concat(
output [4:0] y,
input [2:0]a,b,c
    );
assign y = {a, b[0], c[1]};
endmodule
