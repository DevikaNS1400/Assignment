`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module saturating_add(
input [3:0]a,b,
output [3:0]Y
    );
 wire [4:0]Z ;  
assign Z=a+b;
assign Y=(Z[4])?4'b1111:Z[3:0];
endmodule
