`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
//////////////////////////////////////////////////////////////////////////////////
module mux4_1_tb;
reg [1:0]S;
reg A0,A1,A2,A3;
wire Y;
mux4_1 u1(.Y(Y),.S(S),.A0(A0),.A1(A1),.A2(A2),.A3(A3));
initial begin
$dumpfile("mux4_1_tb.vcd");
$dumpvars(1);
end
initial begin
S=2'b00;A0=1;A1=0;A2=0;A3=0;#10;
S=2'b01;A0=0;A1=1;A2=0;A3=0;#10;
S=2'b10;A0=0;A1=0;A2=1;A3=0;#10;
S=2'b11;A0=0;A1=0;A2=0;A3=1;#10;
$finish;
end
endmodule
