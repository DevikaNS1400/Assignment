`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mux_2_1_tb;
reg I1,I0,S;
wire Y;
mux_2_1_ u1(.Y(Y),.S(S),.I1(I1),.I0(I0));

initial begin
S=0;I1=0;I0=1;#10;
S=1;I1=1;I0=0;#10;
S=0;I1=1;I0=0;#10;
S=1;I1=0;I0=1;#10;
$finish;
end
endmodule
