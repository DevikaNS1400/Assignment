`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module cmos_rpsn_2(
output Y,
input A,B
    );
wire w;
supply0 gnd;
supply1 Vcc;
 pmos p1(w,Vcc,A);
 pmos p2(Y,w,B);
 
 nmos n1(Y,gnd,A);
 nmos n2(Y,gnd,B);
endmodule
