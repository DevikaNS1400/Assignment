`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mux8_1_tb;
reg I0,I1,I2,I3,I4,I5,I6,I7;
reg [2:0]S;
wire Y;
mux_8_1 u4(.Y(Y),.I0(I0),.I1(I1),.I2(I2),.I3(I3),.I4(I4),.I5(I5),.I6(I6),.I7(I7),.S(S));
initial begin
$dumpfile("mux8_1_tb.vcd");
$dumpvars(1);
end
initial 
begin
S=000;I0=1;I1=0;I2=0;I3=0;I4=0;I5=0;I6=0 ;I7=0;#10;
S=001;I0=0;I1=0;I2=0;I3=0;I4=0;I5=0;I6=0;I7=0;#10;
S=010;I0=0;I1=0;I2=1;I3=0;I4=0;I5=0;I6=0;I7=0;#10;
S=011;I0=1;I1=1;I2=0;I3=0;I4=0;I5=0;I6=1;I7=0;#10;
S=100;I0=1;I1=1;I2=0;I3=1;I4=1;I5=0;I6=1;I7=0;#10;
S=101;I0=1;I1=1;I2=0;I3=1;I4=0;I5=0;I6=1;I7=0;#10;
S=110;I0=1;I1=1;I2=0;I3=1;I4=0;I5=0;I6=1;I7=0;#10;
S=111;I0=1;I1=1;I2=0;I3=1;I4=0;I5=0;I6=1;I7=0;#10;
$finish;
end
endmodule