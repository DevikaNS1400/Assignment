`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module zero_one(
output zero,one,
input [7:0]x
    );
    assign zero = ~(|x); 
    assign one = &x;
endmodule
