`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module encoder_4_2_tb;
reg Y3,Y2,Y1,Y0;
wire [1:0]I;
encoder_4_2 u1(.I(I),.Y3(Y3),.Y2(Y2),.Y1(Y1),.Y0(Y0));
initial begin
Y3=0;Y2=0;Y1=1;Y0=0;#10;
Y3=0;Y2=0;Y1=0;Y0=1;#10;
Y3=1;Y2=0;Y1=0;Y0=0;#10;
Y3=0;Y2=1;Y1=0;Y0=0;#10;
Y3=1;Y2=0;Y1=1;Y0=0;#10;
Y3=0;Y2=0;Y1=0;Y0=0;#10;
$finish;
end
endmodule
