`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module buffer_delay(
output y,
input a
);
buf #(3:4:5) g1(y,a);

endmodule
