`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module reg_wire;
reg_module u1();
wire_module u2();
initial
begin
#20;
$finish;
end
endmodule
