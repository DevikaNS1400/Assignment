`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module real_delta_tb;
real_delta u1();
initial begin
$dumpfile("real_delta_tb");
$dumpvars(1);
end
initial begin
#50;
$finish;
end
endmodule
