`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_sum_tb;
wire [3:0]sum;
reg [2:0]a,b;
mod_sum u1(.sum(sum),.a(a),.b(b));
initial begin
a=3'b010;b=3'b101;#10;
a=3'b011;b=3'b111;#10;
a=3'b100;b=3'b111;#10;
a=3'b111;b=3'b101;#10;
$finish;
end
endmodule
