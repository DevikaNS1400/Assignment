`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module parity_gen_tb;
reg [8:0]x;
wire ep,op;
mod_parity u1(.x(x),.ep(ep),.op(op));
initial begin
x=9'b001100110;#10;
x=9'b001110110;#10;
x=9'b101110110;#10;
x=9'b001110110;#10;
$finish;
end
endmodule
