`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_memory();
reg [7:0]mem[0:15];
integer i;
initial begin
i=0;
repeat(16)begin
mem[i]=8'h55;
i=i+1;
end
for (i = 0; i < 16; i = i + 1)
$display("mem[%0d] = %h", i, mem[i]);
end
endmodule