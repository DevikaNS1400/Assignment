`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module cmos_invtr(
output Y,
input A);
supply1 Vcc;
supply0 gnd;

 pmos p1(Y,Vcc,A);
 nmos n1(Y,gnd,A);
endmodule
