`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_operator(
output X,Y,
input [3:0]a,b
    );
assign X=(a==b);
assign Y=(a===b);
endmodule
