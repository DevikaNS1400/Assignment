`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module encoder_4_2(
output [1:0]I,
input Y0,Y1,Y2,Y3
    );
 wire [3:0]c={Y3,Y2,Y1,Y0};  
 assign I=(c==4'b0001)?2'b00:
   (c==4'b0010)?2'b01:
   (c==4'b0100)?2'b10:
   (c==4'b1000)?2'b11:2'bz;
 //assign I=(Y0)?(2'b00):((Y1)?2'b01:((Y2)?2'b10:((Y3)?2'b11:2'bz)));
endmodule
