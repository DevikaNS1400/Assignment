`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module cmos_design1(
output OUT,
input A,B
    );
supply0 gnd;
supply1 Vcc;
wire w1;

pmos p1(OUT,Vcc,A);
pmos p2(OUT,Vcc,B);

nmos n1(w1,gnd,B);
nmos n2(OUT,w1,A);
endmodule
