`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_saturating_tb;
reg [3:0]a,b;
wire [3:0]Y;
saturating_add u1(.Y(Y),.a(a),.b(b));
initial begin
a=4'b0011;b=4'b0111;#10;
a=4'b0111;b=4'b1000;#10;
a=4'b1011;b=4'b0011;#10;
a=4'b1100;b=4'b0100;#10;

$finish;
end
endmodule
