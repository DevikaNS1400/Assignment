`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module bitselect_tb;
bitselect u1();
initial begin
$dumpfile("bitselect_tb.vcd");
$dumpvars(1);
end
initial begin
#30;
end
endmodule
