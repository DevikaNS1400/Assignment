`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_or_operation(
input a,b
    );
assign out = a | b;
endmodule
