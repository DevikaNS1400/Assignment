`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_mux_4_1(
output Y,
input S1,S0,
input i3,i2,i1,i0
    );
 assign Y = S1 ? (S0 ? i3 : i2) : (S0 ? i1 : i0);
endmodule
