`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_sum_tb;
reg [7:0]a,b;
wire [7:0]sum;
mod_tf_sum u1(.sum(sum),.a(a),.b(b));
initial begin
a=3;b=4;#10;
a=6;b=5;#10;
a=2;b=7;#10;
a=10;b=8;#10;
$finish;
end
endmodule
