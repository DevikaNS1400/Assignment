`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_operator_tb;
reg [3:0]a,b;
wire X,Y;
mod_operator u1(.X(X),.Y(Y),.a(a),.b(b));
initial begin
a=4'b10x1;b=4'b10x1;#10;
a=4'b0101;b=4'b1101;#10;
a=4'b1010;b=4'b1010;#10;
a=4'b10z1;b=4'b10z1;#10;
$finish;
end
endmodule
