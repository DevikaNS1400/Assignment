`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_twos_complnt_adr(
output [3:0] sum,
output c_out,
input c_in,
input [3:0]x,y
    );
 wire [3:0] t;
 assign t = y ^ {4{c_in}};
 assign {c_out, sum} = x + t + c_in;   
endmodule
