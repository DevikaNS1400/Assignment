`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_generate_tb;
mod_generate u1();
initial begin 
#30$finish;
end
endmodule
