`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module bitslicing(
output [3:0]W,X,Y,Z,
input [7:0]data);
assign W = data[3:0]+1;
assign X = data[7:4]+1;
assign Y = data[3:0]+4'b0010;
assign Z = data[7:4]+4'b0010;


endmodule
