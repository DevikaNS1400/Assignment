`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
//////////////////////////////////////////////////////////////////////////////////
module mod_demux1_4(
output I3,I2,I1,I0,
input Y,
input [1:0]S,
input en
 );
assign I0 = (en==1&& S==2'b00)?Y:1'b0;
assign I1 = (en==1&& S==2'b01)?Y:1'b0;
assign I2 = (en==1&& S==2'b10)?Y:1'b0;
assign I3 = (en==1&& S==2'b11)?Y:1'b0;
endmodule
