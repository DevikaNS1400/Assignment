
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module comp_tb;
parameter N=4;
reg [N-1:0]a,b;
wire aeb,alb,agb;
mod_N_comp u1(.aeb(aeb),.alb(alb),.agb(agb),.a(a),.b(b));
initial begin
a=1010;b=1101;#10;
a=1010;b=0011;#10;
a=1011;b=1011;#10;
a=1001;b=1100;#10;

$finish;
end
endmodule

