`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mux_2_1_tri(
output Y,
input A,B,S);
bufif0 g1(Y,A,S);
bufif1 g2(Y,B,S);
endmodule
