`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module udp_dlatch_tb;
reg clk,d;
wire q;

udp_d_latch u1(.q(q),.clk(clk),.d(d));

initial begin
clk=0;d=0;#10;
clk=0;d=1;#10;
clk=1;d=0;#10;
clk=1;d=1;#10;
$finish;
end
endmodule
