`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_mux_tb;
reg S1,S0;
reg i3,i2,i1,i0;
wire Y;

mod_mux_4_1 u1(.Y(Y),.S1(S1),.S0(S0),.i3(i3),.i2(i2),.i1(i1),.i0(i0));
initial begin
S1=0;S0=0;i3=0;i2=0;i1=0;i0=1;#10;
S1=0;S0=1;i3=1;i2=1;i1=0;i0=1;#10;
S1=1;S0=0;i3=0;i2=1;i1=0;i0=0;#10;
S1=1;S0=1;i3=0;i2=1;i1=1;i0=1;#10;
$finish;
end
endmodule
