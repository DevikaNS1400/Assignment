`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_n_bit_mux #(parameter N=4)(
output [N-1:0]Y,
input [N-1:0]I0,
input [N-1:0]I1,
input [N-1:0]I2,
input [N-1:0]I3,
input [1:0]S
    );
 assign Y=(S==2'b00)?I0:
          (S==2'b01)?I1:
          (S==2'b10)?I2:
          (S==2'b11)?I3:2'bz;   
endmodule
