`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module decoder_2_4(
input I1,I0,
output y0,y1,y2,y3
    );
 assign y0=I1|I0;
 assign y1=I1|~I0;
 assign y2=~I1|I0;
 assign y3=~I1|~I0;
endmodule
