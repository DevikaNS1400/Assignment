`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_4_bit_fa(
output [3:0]sum,
output c_out,
input [3:0]a,b,
input c_in
    );
assign  {c_out, sum} = a + b + c_in;
endmodule
