`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module priority_encoder_tb;
wire [1:0]S;
reg [3:0]I;
mod_priority_encoder u1(.S(S),.I(I));
initial begin
$monitor("Time=%d I=%b S=%b",$time,I,S);
I=4'b0001;#10;
I=4'b0010;#10;
I=4'b0110;#10;
I=4'b1000;#10;
I=4'b1100;#10;
$finish;
end
endmodule
