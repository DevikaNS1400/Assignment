`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_concat_tb;
reg [2:0]a,b,c;
wire [4:0]y;
mod_concat u1(.y(y),.a(a),.b(b),.c(c));
 initial begin
 a=3'b001;b=3'b110;c=3'b010;#10;
 a=3'b101;b=3'b110;c=3'b111;#10;
 a=3'b001;b=3'b010;c=3'b011;#10;
 a=3'b100;b=3'b101;c=3'b110;#10;
 $finish;
 end
endmodule
