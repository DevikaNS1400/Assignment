`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_shift_left_tb;
wire [7:0]shift_lt;
mod_shift_lt u1(.shift_lt(shift_lt));
initial 
#100$finish;
endmodule
