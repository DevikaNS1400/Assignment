`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module BM_shift_rt_tb;
reg i,clk;
wire y;
bit_shift_reg u1(.y(y),.i(i),.clk(clk));
always 
#5 clk=~clk;
initial
 begin
 clk=0;
 i=0;#10;
 i=1;#10;
 i=1;#10;
 i=0;#10;
 i=1;#10;
 $finish;
 end
endmodule
