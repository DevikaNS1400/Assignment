`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_ab();
reg a,b;  
initial begin a=1; b=a; 
$display($time, "a=%d,b=%d",a,b);  
end  
initial begin #1 a<=1; b<=a;  
$display ($time, "a=%d,b=%d",a,b);  
end  
endmodule
