`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
//////////////////////////////////////////////////////////////////////////////////
module mod_ltrt_shift(
output[3:0] lt_shift_x,rt_shift_x,
input [3:0]x
    );
assign lt_shift_x=(x<<2);
assign rt_shift_x=(x>>2);
endmodule
