`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_nbitmux_tb;
parameter N=4;
reg [N-1:0]I0;
reg [N-1:0]I1;
reg [N-1:0]I2;
reg [N-1:0]I3;
reg [1:0]S;
wire [N-1:0]Y;
mod_n_bit_mux u1(.Y(Y),.I0(I0),.I1(I1),.I2(I2),.I3(I3),.S(S));
initial begin
S=00;I0=4'b0101;I1=4'b1010;I2=4'b0010;I3=0110;#10;
S=01;I0=4'b0101;I1=4'b1010;I2=4'b0010;I3=0110;#10;
S=10;I0=4'b0101;I1=4'b1010;I2=4'b0010;I3=0110;#10;
S=11;I0=4'b0101;I1=4'b1010;I2=4'b0010;I3=0110;#10;
$finish;
end
endmodule
