`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module module_sum(
output sum,
input a,b
    );
assign #5 sum = a + b;

endmodule
