`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_mux_4_1_tb;
reg Y,en;
reg [1:0]S;
wire I3,I2,I1,I0;
mod_demux1_4 u1(.I3(I3),.I2(I2),.I1(I1),.I0(I0),.Y(Y),.en(en),.S(S));
initial begin
en=1'b0;S=2'b00;Y=1'b1;#10;
en=1'b1;S=2'b00;Y=1'b1;#10;
en=1'b1;S=2'b01;Y=1'b1;#10;
en=1'b1;S=2'b10;Y=1'b1;#10;
en=1'b1;S=2'b11;Y=1'b1;#10;
en=1'b0;#10;//S=2'b10;Y=1'b1;#10;
$finish;
end
endmodule
