`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module zero_one_tb;
reg [7:0]x;
wire zero,one;
zero_one u1(.x(x),.zero(zero),.one(one));
initial begin
x=8'b00110011;#10;
x=8'b00000000;#10;
x=8'b10101010;#10;
x=8'b11111111;#10;
$finish;
end
endmodule
