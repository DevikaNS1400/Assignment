`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module register_display_tb;
register_display u1();
initial begin
#20;
end
endmodule
