`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
//////////////////////////////////////////////////////////////////////////////////
module nand_ar_tb;
reg [3:0]a,b;
wire [3:0]nand_ar;

NAND_array u1(.nand_ar(nand_ar),.a(a),.b(b));
initial begin
  $dumpfile("Assignment_1_1Q24_tb.vcd");
  $dumpvars(1);
end
initial begin
a=4'b0110;b=4'b0101;#10;
a=4'b1110;b=4'b1001;#10;
a=4'b0101;b=4'b1011;#10;
a=4'b0111;b=4'b0001;#10;
$finish;
end
endmodule
