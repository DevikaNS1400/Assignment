`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_flag_tb;
reg f1,f2,f3;
wire [2:0]y;
mod_flag u1(.y(y),.f1(f1),.f2(f2),.f3(f3));
initial begin
f3=0;f2=1;f1=1;#10;
f3=1;f2=1;f1=1;#10;
f3=0;f2=1;f1=0;#10;
f3=1;f2=0;f1=0;#10;
f3=1;f2=0;f1=1;#10;
$finish;
end
endmodule
