`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_not(
output y,
input a
    );
    
not #(3,5) g1(y,a)  ;

endmodule
