`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module busmodify_tb;
busmodify u1();
initial begin
$dumpfile("busmodify.vcd");
$dumpvars(1);
end
initial begin
#40;
$finish;
end
endmodule
