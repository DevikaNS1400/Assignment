`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module module_and(
output out,
input a,b  );
assign out=a&b;
endmodule
