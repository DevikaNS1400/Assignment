`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module signed_int_tb;
signed_integer u1();
initial begin
#20;
end
endmodule
