`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_a_b();
reg a,b;
initial begin
a=0;b=0;
end
always@(a,b) begin
//$monitor($time,"a=%d,b=%d",a,b);
#10 a = 1'b0;
#1 b = 1'b1;
a = 1;
#5 b = a;
$display($time,"a=%d,b=%d",a,b);
end
endmodule


/*OUTPUT

16a=1,b=1

*/