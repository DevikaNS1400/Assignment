`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module time_sim_tb;
time_sim u1();
initial begin
#100;
$finish;
end
endmodule
