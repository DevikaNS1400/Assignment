`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module Decoder2_4_tb;
reg I1,I0;
wire y3,y2,y1,y0;
decoder_2_4 u1(.y3(y3),.y2(y2),.y1(y1),.y0(y0),.I1(I1),.I0(I0));
initial
begin
I1=0;I0=0;#10;
I1=0;I0=1;#10;
I1=1;I0=0;#10;
I1=1;I0=1;#10;
$finish;
end
endmodule