`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_dnv_tb;
reg [2:0]a,b;
wire [5:0]m,d;
mod_2function u1(.m(m),.d(d),.a(a),.b(b));
initial begin
a=3'b101;b=3'b011;#10;
a=3'b100;b=3'b111;#10;
a=3'b110;b=3'b010;#10;
a=3'b000;b=3'b001;#10;
$finish;
end
endmodule
