`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_parity(
input [8:0]x,
output ep,op 
    );    
assign ep = ^x;
 assign op = ~ep;
endmodule
