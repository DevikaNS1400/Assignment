`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module register_display();
reg [7:0]A;

initial begin
$display("A=%b",A);
A=01010001;
end
endmodule
