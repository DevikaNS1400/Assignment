`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////

module mod_replication(
output [7:0] y,
input [2:0]a,b,c
    );
assign y = {a, {4{b[0]}}, c[1]};
endmodule
 
