`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module signed_integer();
integer i;
initial begin
i=30;
$display("i=%b",i);
#10;
i=-30;
$display("i=%b",i);
#10;
$finish;
end
endmodule
