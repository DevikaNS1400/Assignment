`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_bitwise(
output [3:0]a,b,c,d,e,
input [3:0]x,y
    );
 assign a=~x;
 assign b=x&y;
 assign c=(x|y);
 assign d=x^y;
 assign e=x^~y;
endmodule
