
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module realtime_sim_tb;
realtime_sim u1();
initial begin
$dumpfile("realtime_sim_tb");
$dumpvars();
end
initial begin
#50;
$finish;
end
endmodule