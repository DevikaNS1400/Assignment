`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_comp(
output ceq,clt,cgt,
input [1:0]C,T
    );
assign ceq=(C==T)?1'b1:1'b0;
assign clt=(C<T)?1'b1:1'b0;
assign cgt=(C>T)?1'b1:1'b0;
endmodule
