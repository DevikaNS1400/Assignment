`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_mem_tb;
mod_memory u1();
initial begin
#40$finish;
end
endmodule
