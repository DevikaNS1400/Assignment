`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module part_select_tb;
part_select u1();
initial begin
$dumpfile("part_select_tb.vcd");
$dumpvars(1);
end
initial begin
#40;
$finish;
end
endmodule
