`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_clk(
    );
reg clk;
initial clk=0;
initial begin
forever #5 clk=~clk;
end
endmodule
