`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module part_select();
reg [7:0]bus;
initial begin
bus=8'b01011101;
$display("The lower nibble bus[3:0]=%b",bus[3:0]);#10;
$finish;
end
endmodule
