`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_casex_tb;
reg I0,I1,I2,I3,I4,I5,I6,I7;
reg [2:0]s;
wire y;
mod_casex u1(.y(y),.s(s),.I0(I0),.I1(I1),.I2(I2),.I3(I3),.I4(I4),.I5(I5),.I6(I6),.I7(I7));
initial begin
s=000;I0=1;I1=0;I2=0;I3=0;I4=0;I5=0;I6=0;I7=0;#10;
s=001;I0=0;I1=1;I2=0;I3=0;I4=0;I5=0;I6=0;I7=0;#10;
s=010;I0=0;I1=0;I2=1;I3=0;I4=0;I5=0;I6=0;I7=0;#10;
s=011;I0=0;I1=0;I2=0;I3=1;I4=0;I5=0;I6=0;I7=0;#10;
s=100;I0=0;I1=0;I2=0;I3=0;I4=1;I5=0;I6=0;I7=0;#10;
s=101;I0=0;I1=0;I2=0;I3=0;I4=0;I5=1;I6=0;I7=0;#10;
s=110;I0=0;I1=0;I2=0;I3=0;I4=0;I5=0;I6=1;I7=0;#10;
s=111;I0=0;I1=0;I2=0;I3=0;I4=0;I5=0;I6=0;I7=1;#10;
$finish;
end
endmodule
