`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mux_4_1_tb;
reg I3,I2,I1,I0,S1,S0;
wire Y;

mux_4_1 u1(.Y(Y),.S1(S1),.S0(S0),.I3(I3),.I2(I2),.I1(I1),.I0(I0));
initial begin
S1=0;S0=0;I3=1;I2=1;I1=1;I0=0;#10;
S1=0;S0=1;I3=0;I2=0;I1=1;I0=0;#10;
S1=1;S0=0;I3=1;I2=0;I1=1;I0=1;#10;
S1=1;S0=1;I3=1;I2=0;I1=0;I0=0;#10;
$finish;
end
endmodule
