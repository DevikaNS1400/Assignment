`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_comp_tb;
reg [1:0]C,T;
wire ceq,clt,cgt;
mod_comp u1(.ceq(ceq),.clt(clt),.cgt(cgt),.C(C),.T(T));
initial begin
C=10;T=00;#10;
C=11;T=11;#10;
C=01;T=10;#10;
C=10;T=10;#10;
$finish;
end
endmodule
