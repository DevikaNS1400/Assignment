`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module bitselect();
reg [7:0]data;

initial begin
data=8'b10101100;
$display("The value at data[3]=%b",data[3]);
end

endmodule
