`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module cmos_invtr_tb;
reg A;
wire Y;
cmos_invtr u1(.Y(Y),.A(A));
initial begin
$dumpfile("cmos_invtr_tb.vcd");
$dumpvars(1);
end
initial begin
A=0;#10;
A=1;#10;
$finish;
end
endmodule
