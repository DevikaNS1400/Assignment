`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mux_2_1_(
output Y,
input I1,I0,
input S
    );
    
assign Y= (S)?I1:I0;
endmodule
