`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module mod_shift_rt_tb;
reg [4:0]x;
wire [4:0]y;
mod_f_shiftrt u1(.y(y),.x(x));
initial begin
x=5'b0100;#10;
x=5'b1000;#10;
x=5'b0010;#10;
x=5'b0001;#10;
$finish;
end
endmodule
